

library  IEEE;
use      IEEE.std_logic_1164.all;
use 	 IEEE.STD_LOGIC_UNSIGNED.ALL;
use 	 ieee.numeric_std.all;



entity transmit_arp_reply is
   port (clk_i :         in   std_logic;
         start_i :       in   std_logic;
         reset_i :       in   std_logic;
		 MAC_src_addr_i :  in   std_logic_vector(47 downto 0);
		 tell_MAC_addr_i :  in   std_logic_vector(47 downto 0);
		 IP_src_addr_i :  in   std_logic_vector(31 downto 0);
		 tell_IPaddr_i :  in   std_logic_vector(31 downto 0);
		
         ff_tx_data_o :         out  std_logic_vector(7 downto 0);  
         ff_tx_valid_o :        out  std_logic;
         ff_tx_last_o :         out  std_logic);
 		
end transmit_arp_reply;



architecture rtl of transmit_arp_reply is


  type t_state is (waiting,
                   H_01, H_02, H_03, H_04,
                   H_11, H_12, H_13, H_14,
                   H_21, H_22, H_23, H_24,
                   H_31, H_32, H_33, H_34,
                   H_41, H_42, H_43, H_44,
                   H_51, H_52, H_53, H_54,
                   H_61, H_62, H_63, H_64,
                   H_71, H_72, H_73, H_74,
                   H_81, H_82, H_83, H_84,
                   H_91, H_92, H_93, H_94,
                   H_101, H_102, H_103, H_104,
                   
				   payload_11, payload_12, payload_13, payload_14,
				   payload_21, payload_22, payload_23, payload_24,
				   payload_31, payload_32, payload_33, payload_34,
				   payload_41, payload_42, payload_43, payload_44,
                   eop1, eop2, eop3, eop4,
                   terminate);
		
		
  signal s_state : t_state;
  signal s_ff_tx_wren_o :std_logic;
 
  
begin    

 
  
p_ctrl: process (clk_i, reset_i)
begin  -- process p_serin
  if (reset_i = '1') then               -- asynchronous reset (active high)
    s_state <= waiting;
    ff_tx_data_o <=  x"00";
    ff_tx_data_o <=  x"00";
    ff_tx_last_o <= '0';
    s_ff_tx_wren_o <= '0';
   
  elsif rising_edge(clk_i) then  -- rising clock edge
    case s_state is
    
        when H_01 =>    ff_tx_data_o <= tell_MAC_addr_i(47 downto 40);  s_ff_tx_wren_o <= '1';  s_state <= H_02;
        when H_02 =>    ff_tx_data_o <= tell_MAC_addr_i(39 downto 32); 		                    s_state <= H_11;
            
	    when H_11 =>	ff_tx_data_o <=  tell_MAC_addr_i(31 downto 24);					        s_state <= H_12;
	    when H_12 =>	ff_tx_data_o <=  tell_MAC_addr_i(23 downto 16);					        s_state <= H_13;
	    when H_13 =>	ff_tx_data_o <=  tell_MAC_addr_i(15 downto 8);					        s_state <= H_14;
	    when H_14 =>	ff_tx_data_o <=  tell_MAC_addr_i(7 downto 0);					        s_state <= H_21;
	    
		when H_21 =>    ff_tx_data_o <=  MAC_src_addr_i(47 downto 40);							s_state <= H_22;
		when H_22 =>    ff_tx_data_o <=  MAC_src_addr_i(39 downto 32);							s_state <= H_23;
		when H_23 =>    ff_tx_data_o <=  MAC_src_addr_i(31 downto 24);							s_state <= H_24;
		when H_24 =>    ff_tx_data_o <=  MAC_src_addr_i(23 downto 16);							s_state <= H_31;
		
		when H_31 =>	ff_tx_data_o <=  MAC_src_addr_i(15 downto 8);                           s_state <= H_32; 
		when H_32 =>	ff_tx_data_o <=  MAC_src_addr_i(7 downto 0);                            s_state <= H_33; 
		when H_33 =>	ff_tx_data_o <=  x"08";                                                 s_state <= H_34; 
		when H_34 =>	ff_tx_data_o <=  x"06";                                                 s_state <= H_41;
		
		when H_41 =>    ff_tx_data_o <=  x"00"; 					            	            s_state <= H_42;
		when H_42 =>    ff_tx_data_o <=  x"01";						                            s_state <= H_43;
		when H_43 =>    ff_tx_data_o <=  x"08";	                        				        s_state <= H_44;
		when H_44 =>    ff_tx_data_o <=  x"00"; 		                				        s_state <= H_51;
		
		when H_51 =>	ff_tx_data_o <=  x"06";				                                  	s_state <= H_52;
		when H_52 =>	ff_tx_data_o <=  x"04";				                                    s_state <= H_53;
		when H_53 =>	ff_tx_data_o <=  x"00";			                                        s_state <= H_54;
		when H_54 =>	ff_tx_data_o <=  x"02";				                          			s_state <= H_61;
		
		when H_61 =>    ff_tx_data_o <=  MAC_src_addr_i(47 downto 40);							s_state <= H_62;
		when H_62 =>    ff_tx_data_o <=  MAC_src_addr_i(39 downto 32);							s_state <= H_63;
		when H_63 =>    ff_tx_data_o <=  MAC_src_addr_i(31 downto 24);							s_state <= H_64;
		when H_64 =>    ff_tx_data_o <=  MAC_src_addr_i(23 downto 16);							s_state <= H_71;
		
		when H_71 =>	ff_tx_data_o <=  MAC_src_addr_i(15 downto 8);                           s_state <= H_72; 
		when H_72 =>	ff_tx_data_o <=  MAC_src_addr_i(7 downto 0);                            s_state <= H_73; 
		when H_73 =>	ff_tx_data_o <=  IP_src_addr_i(31 downto 24);                           s_state <= H_74; 
		when H_74 =>	ff_tx_data_o <=  IP_src_addr_i(23 downto 16);                           s_state <= H_81;
		
		when H_81 =>	ff_tx_data_o <=  IP_src_addr_i(15 downto 8);			 				s_state <= H_82;
		when H_82 =>	ff_tx_data_o <=  IP_src_addr_i(7 downto 0);			  	    			s_state <= H_83;
		when H_83 =>	ff_tx_data_o <=  tell_MAC_addr_i(47 downto 40);			  				s_state <= H_84;
		when H_84 =>	ff_tx_data_o <=  tell_MAC_addr_i(39 downto 32);                         s_state <= H_91;
		
		when H_91 =>	ff_tx_data_o <=  tell_MAC_addr_i(31 downto 24);					        s_state <= H_92;
	    when H_92 =>	ff_tx_data_o <=  tell_MAC_addr_i(23 downto 16);					        s_state <= H_93;
	    when H_93 =>	ff_tx_data_o <=  tell_MAC_addr_i(15 downto 8);					        s_state <= H_94;
	    when H_94 =>	ff_tx_data_o <=  tell_MAC_addr_i(7 downto 0);					        s_state <= H_101;
	    
	    when H_101 =>	ff_tx_data_o <=  tell_IPaddr_i(31 downto 24);					        s_state <= H_102;
	    when H_102 =>	ff_tx_data_o <=  tell_IPaddr_i(23 downto 16);					        s_state <= H_103;
	    when H_103 =>	ff_tx_data_o <=  tell_IPaddr_i(15 downto 8);					        s_state <= H_104;
	    when H_104 =>	ff_tx_data_o <=  tell_IPaddr_i(7 downto 0);					            s_state <= payload_11;
      
		when payload_11 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_12;
		when payload_12 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_13;
		when payload_13 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_14;
		when payload_14 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_21;
		
		when payload_21 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_22;
		when payload_22 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_23;
		when payload_23 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_24;
		when payload_24 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_31;
		
		when payload_31 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_32;
		when payload_32 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_33;
		when payload_33 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_34;
		when payload_34 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_41;
		
		when payload_41 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_42;
		when payload_42 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_43;
		when payload_43 =>		ff_tx_data_o <=  x"00";         								s_state <= payload_44;
		when payload_44 =>		ff_tx_data_o <=  x"00";         								s_state <= eop3;
		
--		when eop1 =>	    	ff_tx_data_o <=  x"00";         								s_state <= eop2;
--		when eop2 =>	    	ff_tx_data_o <=  x"00";         								s_state <= eop3;
		when eop3 =>	    	ff_tx_data_o <=  x"00";         								s_state <= eop4;
		when eop4 =>		    ff_tx_data_o <=  x"00";    ff_tx_last_o <= '1';					s_state <= terminate;	
      ---------------------------------------------------------------------------------------------------------------------------------------------------
		when terminate =>	ff_tx_data_o <=  x"00";	 s_ff_tx_wren_o <= '0';	ff_tx_last_o <='0'; s_state <= waiting ;
      ---------------------------------------------------------------------------------------------------------------------------------------------------
      
      
      when others =>
        if start_i = '1' then
          -- START Condition detected
          s_state <= H_01;
          
        end if;
    end case;
  end if;
end process p_ctrl;

ff_tx_valid_o <= s_ff_tx_wren_o;

end rtl;
